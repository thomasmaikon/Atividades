module xore(x1,x2,saida);
		
		input logic x1,x2;
		output logic saida;
		
		assign saida = x1 ^ x2;
		
endmodule
